* Extracted by KLayout with SG13G2 LVS runset on : 04/07/2025 15:23

.SUBCKT tg_layout_v2
X$1 \$3 \$4 \$3 \$4 \$1 nmos
X$2 \$3 \$4 \$3 \$2 \$1 pmos$1
.ENDS tg_layout_v2

.SUBCKT pmos$1 \$3 \$4 \$5 \$8 \$9
M$1 \$2 \$1 \$3 \$8 sg13_lv_pmos L=0.13u W=10u AS=3.4p AD=1.9p PS=20.68u
+ PD=10.38u
M$2 \$3 \$7 \$4 \$8 sg13_lv_pmos L=0.13u W=10u AS=1.9p AD=1.9p PS=10.38u
+ PD=10.38u
M$3 \$4 \$10 \$5 \$8 sg13_lv_pmos L=0.13u W=10u AS=1.9p AD=3.4p PS=10.38u
+ PD=20.68u
.ENDS pmos$1

.SUBCKT nmos \$1 \$2 \$3 \$4 \$5
M$1 \$1 \$7 \$2 \$5 sg13_lv_nmos L=0.13u W=4u AS=1.36p AD=0.76p PS=8.68u
+ PD=4.38u
M$2 \$2 \$8 \$3 \$5 sg13_lv_nmos L=0.13u W=4u AS=0.76p AD=0.76p PS=4.38u
+ PD=4.38u
M$3 \$3 \$9 \$4 \$5 sg13_lv_nmos L=0.13u W=4u AS=0.76p AD=1.36p PS=4.38u
+ PD=8.68u
.ENDS nmos
